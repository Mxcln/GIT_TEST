module mod_yyd(
    input a,
    output b
);
    assign b =a;
endmodule