#module  #(
    parameters
) (
    ports
);
    
endmodule